
module peripheral_control_movimiento_TB;

  
  
  
   reg clk;
   reg rst;
   reg [15:0]d_in;
   reg cs;
   reg [3:0]addr;
   reg rd;
   reg wr;
   wire [15:0]d_out;



  peripheral_control_movimiento  uut (.clk(clk), 
				         .rst(rst), 
					 .d_in(d_in), 
					 .cs(cs), 
					 .addr(addr), 
					 .rd(rd), 
					 .wr(wr), 
					 .d_out(d_out));

//inicialización 


parameter PERIOD          = 20;
parameter real DUTY_CYCLE = 0.5;
parameter OFFSET          = 0;
reg [20:0] i;
event reset_trigger;


   initial begin  // Initialize Inputs
      clk = 0; rst = 1; d_in = 16'd0035; addr = 16'h0000; cs=1; rd=0; wr=1; 
   end


 initial  begin  // Process for clk
     #OFFSET;
     forever
       begin
         clk = 1'b0;
         #(PERIOD-(PERIOD*DUTY_CYCLE)) clk = 1'b1;
         #(PERIOD*DUTY_CYCLE);
       end
   end




   initial begin: TEST_CASE
     $dumpfile("peripheral_control_movimiento_TB.vcd");
    $dumpvars(-1, uut);
	
     #10 -> reset_trigger;
     #((PERIOD*DUTY_CYCLE)*200) $finish;
   end

endmodule
